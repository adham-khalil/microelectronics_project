part_a.end

.include MOSFET_models_0p5_0p18-1.inc

VIN vi gnd PULSE(0 1.8 0.5n 1p 1p 20n)
VDD vdd gnd DC 1.8
* Transistors
M1 vo vi gnd gnd NMOS0P18 [w=0.9u l=0.18u]
M2 vo vi vdd vdd PMOS0P18 [w=0.9u l=0.18u]

* Load
RL vo vc 1k
CL vc gnd .2p

.tran 5n 40n
.op
