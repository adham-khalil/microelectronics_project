part_a_matched.end

.include MOSFET_models_0p5_0p18-1.inc

VIN vi gnd 0
VDD vdd gnd DC 1.8
* Transistors
M1 vo vi gnd gnd NMOS0P18 [w=0.9u l=0.18u]
M2 vo vi vdd vdd PMOS0P18 [w=2.25u l=0.18u]

* Load
RL vo vc 1k
CL vc gnd .2p

* DC Sweep Analysis
.dc VIN 0 1.8 0.01
.op
